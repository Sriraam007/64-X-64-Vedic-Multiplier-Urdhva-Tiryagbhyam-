module Full_Adder_64bit(A,B,cin,SUM,cout);
    input [63:0]A,B;
    input cin;
    output [63:0]SUM;
    output cout;
    wire [63:0]w;
    
    Full_Adder2 F1(A[0],B[0],cin,SUM[0],w[0]);
    Full_Adder2 F2(A[1],B[1],w[0],SUM[1],w[1]);
    Full_Adder2 F3(A[2],B[2],w[1],SUM[2],w[2]);
    Full_Adder2 F4(A[3],B[3],w[2],SUM[3],w[3]);
    Full_Adder2 F5(A[4],B[4],w[3],SUM[4],w[4]);
    Full_Adder2 F6(A[5],B[5],w[4],SUM[5],w[5]);
    Full_Adder2 F7(A[6],B[6],w[5],SUM[6],w[6]);
    Full_Adder2 F8(A[7],B[7],w[6],SUM[7],w[7]);
    Full_Adder2 F9(A[8],B[8],w[7],SUM[8],w[8]);
    Full_Adder2 F10(A[9],B[9],w[8],SUM[9],w[9]);
    Full_Adder2 F11(A[10],B[10],w[9],SUM[10],w[10]);
    Full_Adder2 F12(A[11],B[11],w[10],SUM[11],w[11]);
    Full_Adder2 F13(A[12],B[12],w[11],SUM[12],w[12]);
    Full_Adder2 F14(A[13],B[13],w[12],SUM[13],w[13]);
    Full_Adder2 F15(A[14],B[14],w[13],SUM[14],w[14]);
    Full_Adder2 F16(A[15],B[15],w[14],SUM[15],w[15]);
    
    Full_Adder2 F17(A[16],B[16],w[15],SUM[16],w[16]);
    Full_Adder2 F18(A[17],B[17],w[16],SUM[17],w[17]);
    Full_Adder2 F19(A[18],B[18],w[17],SUM[18],w[18]);
    Full_Adder2 F20(A[19],B[19],w[18],SUM[19],w[19]);
    Full_Adder2 F21(A[20],B[20],w[19],SUM[20],w[20]);
    Full_Adder2 F22(A[21],B[21],w[20],SUM[21],w[21]);
    Full_Adder2 F23(A[22],B[22],w[21],SUM[22],w[22]);
    Full_Adder2 F24(A[23],B[23],w[22],SUM[23],w[23]);
    Full_Adder2 F25(A[24],B[24],w[23],SUM[24],w[24]);
    Full_Adder2 F26(A[25],B[25],w[24],SUM[25],w[25]);
    Full_Adder2 F27(A[26],B[26],w[25],SUM[26],w[26]);
    Full_Adder2 F28(A[27],B[27],w[26],SUM[27],w[27]);
    Full_Adder2 F29(A[28],B[28],w[27],SUM[28],w[28]);
    Full_Adder2 F30(A[29],B[29],w[28],SUM[29],w[29]);
    Full_Adder2 F31(A[30],B[30],w[29],SUM[30],w[30]);
    Full_Adder2 F32(A[31],B[31],w[30],SUM[31],w[31]);
    
    Full_Adder2 F33(A[32],B[32],w[31],SUM[32],w[32]);
    Full_Adder2 F34(A[33],B[33],w[32],SUM[33],w[33]);
    Full_Adder2 F35(A[34],B[34],w[33],SUM[34],w[34]);
    Full_Adder2 F36(A[35],B[35],w[34],SUM[35],w[35]);
    Full_Adder2 F37(A[36],B[36],w[35],SUM[36],w[36]);
    Full_Adder2 F38(A[37],B[37],w[36],SUM[37],w[37]);
    Full_Adder2 F39(A[38],B[38],w[37],SUM[38],w[38]);
    Full_Adder2 F40(A[39],B[39],w[38],SUM[39],w[39]);
    Full_Adder2 F41(A[40],B[40],w[39],SUM[40],w[40]);
    Full_Adder2 F42(A[41],B[41],w[40],SUM[41],w[41]);
    Full_Adder2 F43(A[42],B[42],w[41],SUM[42],w[42]);
    Full_Adder2 F44(A[43],B[43],w[42],SUM[43],w[43]);
    Full_Adder2 F45(A[44],B[44],w[43],SUM[44],w[44]);
    Full_Adder2 F46(A[45],B[45],w[44],SUM[45],w[45]);
    Full_Adder2 F47(A[46],B[46],w[45],SUM[46],w[46]);
    Full_Adder2 F48(A[47],B[47],w[46],SUM[47],w[47]);
    
    Full_Adder2 F49(A[48],B[48],w[47],SUM[48],w[48]);
    Full_Adder2 F50(A[49],B[49],w[48],SUM[49],w[49]);
    Full_Adder2 F51(A[50],B[50],w[49],SUM[50],w[50]);
    Full_Adder2 F52(A[51],B[51],w[50],SUM[51],w[51]);
    Full_Adder2 F53(A[52],B[52],w[51],SUM[52],w[52]);
    Full_Adder2 F54(A[53],B[53],w[52],SUM[53],w[53]);
    Full_Adder2 F55(A[54],B[54],w[53],SUM[54],w[54]);
    Full_Adder2 F56(A[55],B[55],w[54],SUM[55],w[55]);
    Full_Adder2 F57(A[56],B[56],w[55],SUM[56],w[56]);
    Full_Adder2 F58(A[57],B[57],w[56],SUM[57],w[57]);
    Full_Adder2 F59(A[58],B[58],w[57],SUM[58],w[58]);
    Full_Adder2 F60(A[59],B[59],w[58],SUM[59],w[59]);
    Full_Adder2 F61(A[60],B[60],w[59],SUM[60],w[60]);
    Full_Adder2 F62(A[61],B[61],w[60],SUM[61],w[61]);
    Full_Adder2 F63(A[62],B[62],w[61],SUM[62],w[62]);
    Full_Adder2 F64(A[63],B[63],w[62],SUM[63],w[63]);
    
    
    assign cout=w[63];
endmodule
